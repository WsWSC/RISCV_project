module top(
    
);




endmodule