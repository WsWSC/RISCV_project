module pc_reg(
    input wire clk,
    input wire rst,

    output reg[31:0] pc_o

);



endmodule