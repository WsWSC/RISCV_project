**************************************************
* risc v side project                            *
*                                                *
* create by WsWSC                                *
**************************************************

module if_id(
    input wire clk,
    input wire rst,
    input wire[31:0] inst_i,
    input wire[31:0] inst_addr_i,

    output wire[31:0] inst_addr_o,
    output wire[31:0] inst_o
);


endmodule