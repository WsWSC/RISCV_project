module dual_ram #(
    parameters;
) (
    input  ;
);
    
endmodule