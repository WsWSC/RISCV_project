**************************************************
* risc v side project                            *
*                                                *
* create by WsWSC                                *
**************************************************

module(

);


endmodule